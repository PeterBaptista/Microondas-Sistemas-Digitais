module encoder( input wire [9:0] keypad,
                input wire enablen,
                input wire clk,
                output wire [3:0] bcd_output,
                input wire load,
                )


endmodule