`include "counter_mod6.v"
`include "counter_mod10.v"

module timer();


endmodule
