module microwave(
    input wire start,
    input wire stopn,
    input wire clearn,
    input wire door_closed,
    input wire [9:0] keypad,
    input wire clk,
    output wire [6:0] second_units_display,
    output wire [6:0] second_tens_display,
    output wire [6:0] minutes_display
)


endmodule